
.include TSMC180.lib

.model pch_tt pmos
.model nch_tt nmos

Vsrc Vdd  0 1.8

.param beta = 6.67

MN1 o1 out 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP1 o1 out Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u

MN2 o2 o1 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP2 o2 o1 Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u

MN3 o3 o2 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP3 o3 o2 Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u

MN4 o4 o3 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP4 o4 o3 Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u

MN5 o5 o4 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP5 o5 o4 Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u

MN6 o6 o5 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP6 o6 o5 Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u

MN7 out o6 0 	0 	nch_tt 	W = 0.18u	L = 0.18u 
MP7 out o6 Vdd 	Vdd	pch_tt	W = beta*0.18u	L = 0.18u




.control


	

tran 1p 5n uic
run 
meas TRAN T_period trig V(out) Val = 1 cross = 3 targ V(out) val = 1 cross = 5

let f = 1/T_period
let tp = T_period/(2*7)
print f

plot V(out)


wrdata 2.a.dat V(out) 
.endc
.end 
