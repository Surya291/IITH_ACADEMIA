* netlist

.include TSMC180.lib


.model nch_tt nmos (level = 8)

Vgs	g	0	2
Vds	d	a	1

V_am	a	0	0

*Ms	d	g	0	0	nch_tt	W=0.27u L=0.18u
Ml	d	g	0	0	nch_tt	W=15u L = 10u

.control


dc Vds 0 1.8  0.005    Vgs 1 2 0.5  

plot -i(V_am) title  "Short Channel"

wrdata 4.1.b.dat -i(V_am)
.endc

.end	



	

