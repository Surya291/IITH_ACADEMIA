*** For Ques: 1
*** NMOS:  W/L = 240/180
*** Vgs = 1.8V, init Vds = 1.8V.,  


.include TSMC180.lib
.model nch_tt nmos (level = 8)

Vgs	g	0	1.8   
V_am	d	am	0V   	** ammeter   
C	am	0	1e-12  	IC = 1.8V 
*R	am	0	1e0
M1	d	g	0	0  nch_tt   W=240n  L = 180n

.ic V(am) = 1.8V
.control

tran 1p  13n 
*plot V(am)
*plot -i(V_am) vs V(am)  title "I vs V"
plot V(am)/-i(V_am) vs V(am) title " Res vs V " 

.endc
.end
