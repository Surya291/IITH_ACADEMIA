***  1st question.. 
***  Varying scaling factor..

.include TSMC180.lib

.model pch_tt pmos
.model nch_tt nmos

*** below for NO-LOAD
Vin inp 0 PULSE( 1.8 3p 3p  3p  3p 500p 1n )
*** below for C-load
*Vin inp 0 PULSE( 1.8 0 0  0  0 1u 2u )
*C out 0  20p

Vsrc  Vdd	0  dc  1.8
MN out inp 0 	0 	nch_tt 	W =0.18u	L = 0.18u 
MP out inp Vdd 	Vdd	pch_tt	W = 0.18u	L = 0.18u


*** While loop to loop over diff values of s and find the prop delay..



.control

let tlhs = vector(20)
let thls = vector(20)
let tps = vector (20)
let s_factor = vector(20)
let loop = 1

while loop < 21 
*** looping 20 times
	let beta = 6
	alter @MN W=loop*0.18u
	alter @MP W=loop*beta*0.18u
	
	*** Uncomment for noload
	tran .1p 5n

	*** Uncomment for load
	*tran  1n 5u
	run

	meas tran O_max max out
	meas tran I_max max inp

	let I_half = 0.5*I_max
	let O_half = 0.5*O_max


	meas tran tplh	trig V(inp) VAL = I_half CROSS=3 targ V(out) VAL=O_half CROSS=3 
	meas tran tphl  trig V(inp) VAL = I_half CROSS=4 targ V(out) VAL=O_half CROSS=4 

	let tp = (tplh + tphl) * 0.5
	
	let tlhs[loop-1] = tplh
	let thls[loop-1] = tphl
	let tps[loop-1] = tp
	let s_factor[loop-1] = loop

	let loop = loop+1
end
plot tps vs s_factor
plot V(out)

*wrdata 1.a.1.dat s_factor vs tps
wrdata 1.a.2.dat s_factor vs tps

.endc
.end










